library verilog;
use verilog.vl_types.all;
entity beat_Cycle_vlg_vec_tst is
end beat_Cycle_vlg_vec_tst;
