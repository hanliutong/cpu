library verilog;
use verilog.vl_types.all;
entity CLK_maker_vlg_check_tst is
    port(
        clk             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end CLK_maker_vlg_check_tst;
