library verilog;
use verilog.vl_types.all;
entity Timer_vlg_vec_tst is
end Timer_vlg_vec_tst;
