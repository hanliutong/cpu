library verilog;
use verilog.vl_types.all;
entity X_IBUS_vlg_vec_tst is
end X_IBUS_vlg_vec_tst;
