module R_addr(
input d,
input [2:0]_reg,
input [2:0]r_m,
input w,DST,EXC,
input [1:0]MOD,
input [3:0]T,
output reg [15:0]R
);
wire Beat,D_E;
assign Beat = T[0]||T[1]||T[2]||T[3];
assign D_E =  DST||EXC;
assign MD = MOD[0]&&MOD[1];

always @ (D_E or Beat or w or d or _reg or r_m or MD)
begin
	if ((D_E&&d)||(!D_E&&!d))
	begin
		case({_reg,w})
		4'b000_0:R=16'b1000000000000000;
		4'b000_1:R=16'b0100000000000000;
		4'b001_0:R=16'b0010000000000000;
		4'b001_1:R=16'b0001000000000000;
		4'b010_0:R=16'b0000100000000000;
		4'b010_1:R=16'b0000010000000000;
		4'b011_0:R=16'b0000001000000000;
		4'b011_1:R=16'b0000000100000000;
		4'b100_0:R=16'b0000000010000000;
		4'b100_1:R=16'b0000000001000000;
		4'b101_0:R=16'b0000000000100000;
		4'b101_1:R=16'b0000000000010000;
		4'b110_0:R=16'b0000000000001000;
		4'b110_1:R=16'b0000000000000100;
		4'b111_0:R=16'b0000000000000010;
		4'b111_1:R=16'b0000000000000001;
		default:R=16'b000000000000000;
		endcase
	end
	else if ((D_E&&!d&&MD)||(!D_E&&d&&MD))
	begin
		case({r_m,w})
		4'b000_0:R=16'b1000000000000000;
		4'b000_1:R=16'b0100000000000000;
		4'b001_0:R=16'b0010000000000000;
		4'b001_1:R=16'b0001000000000000;
		4'b010_0:R=16'b0000100000000000;
		4'b010_1:R=16'b0000010000000000;
		4'b011_0:R=16'b0000001000000000;
		4'b011_1:R=16'b0000000100000000;
		4'b100_0:R=16'b0000000010000000;
		4'b100_1:R=16'b0000000001000000;
		4'b101_0:R=16'b0000000000100000;
		4'b101_1:R=16'b0000000000010000;
		4'b110_0:R=16'b0000000000001000;
		4'b110_1:R=16'b0000000000000100;
		4'b111_0:R=16'b0000000000000010;
		4'b111_1:R=16'b0000000000000001;
		default:R=16'b000000000000000;
		endcase
	end
	else
	begin
		if(Beat)
		begin
			case(r_m)
				3'b000:R=16'b0000000100000000;
				3'b001:R=16'b0000000100000000;
				3'b010:R=16'b0000000000010000;
				3'b011:R=16'b0000000000010000;
				3'b100:R=16'b0000000000000100;
				3'b101:R=16'b0000000000000001;
				3'b110:R=16'b0000000000010000;
				3'b111:R=16'b0000000100000000;
			default:R=16'b000000000000000;
			endcase
		end
		else
		begin
			case(r_m)
				3'b000:R=16'b0000000000000100;
				3'b001:R=16'b0000000000000001;
				3'b010:R=16'b0000000000000100;
				3'b011:R=16'b0000000000000001;
				3'b100:R=16'b0000000000000100;
				3'b101:R=16'b0000000000000001;
				3'b110:R=16'b0000000000010000;
				3'b111:R=16'b0000000100000000;
			default:R=16'b000000000000000;
			endcase
		end
	end

end

endmodule
