module ModRM2R(RM,mod,beat,R);
input [2:0]RM;
input mod,beat;
output reg [15:0]R;
always @ (RM or beat or mod)
if(mod) R=16'b0000000000000000;
else if(beat)
	begin
		case(RM)
			3'b000:R=16'b0000000100000000;
			3'b001:R=16'b0000000100000000;
			3'b010:R=16'b0000000000010000;
			3'b011:R=16'b0000000000010000;
			3'b100:R=16'b0000000000000100;
			3'b101:R=16'b0000000000000001;
			3'b110:R=16'b0000000000010000;
			3'b111:R=16'b0000000100000000;
		default:R=16'b000000000000000;
		endcase
	end
else
		begin
		case(RM)
			3'b000:R=16'b0000000000000100;
			3'b001:R=16'b0000000000000001;
			3'b010:R=16'b0000000000000100;
			3'b011:R=16'b0000000000000001;
			3'b100:R=16'b0000000000000100;
			3'b101:R=16'b0000000000000001;
			3'b110:R=16'b0000000000010000;
			3'b111:R=16'b0000000100000000;
		default:R=16'b000000000000000;
		endcase
	end

endmodule
