library verilog;
use verilog.vl_types.all;
entity R_adrr_vlg_vec_tst is
end R_adrr_vlg_vec_tst;
