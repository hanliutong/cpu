library verilog;
use verilog.vl_types.all;
entity MyCPU is
    port(
        FI              : out    vl_logic;
        DST             : out    vl_logic;
        SRC             : out    vl_logic;
        EXC             : out    vl_logic;
        INT             : out    vl_logic;
        CLK             : out    vl_logic;
        OpCode          : out    vl_logic_vector(5 downto 0);
        IBUS_IR         : out    vl_logic;
        IBUS            : out    vl_logic_vector(15 downto 0);
        ALU_IBUS        : out    vl_logic;
        ADDC            : out    vl_logic;
        SUBC            : out    vl_logic;
        INCAC           : out    vl_logic;
        DECAC           : out    vl_logic;
        W_B             : out    vl_logic;
        IBUS_RA         : out    vl_logic;
        IBUS_RB         : out    vl_logic;
        MDR_DBUS        : out    vl_logic;
        MDR_IBUS        : out    vl_logic;
        BUS_MDR         : out    vl_logic;
        I_DBUS          : out    vl_logic;
        DBUS            : out    vl_logic_vector(15 downto 0);
        MRD             : out    vl_logic;
        MWR             : out    vl_logic;
        M_clk           : out    vl_logic;
        ABUS            : out    vl_logic_vector(15 downto 0);
        MAR_ABUS        : out    vl_logic;
        MAR_IBUS        : out    vl_logic;
        IBUS_MAR        : out    vl_logic;
        IBUS_SR         : out    vl_logic;
        SR_IBUS         : out    vl_logic;
        R_IBUS          : out    vl_logic;
        RE              : out    vl_logic;
        WE              : out    vl_logic;
        R               : out    vl_logic_vector(15 downto 0);
        T               : out    vl_logic_vector(7 downto 0);
        Start           : in     vl_logic;
        IBUS_RBL        : out    vl_logic;
        RBL_IBUS        : out    vl_logic;
        PC_IBUS         : out    vl_logic;
        PCplus1         : out    vl_logic;
        IBUS_PC         : out    vl_logic;
        zero_PC         : out    vl_logic;
        Crystal         : in     vl_logic;
        setTp1          : out    vl_logic;
        A_plus          : out    vl_logic_vector(15 downto 0);
        cnt             : out    vl_logic_vector(3 downto 0);
        jieguo          : out    vl_logic_vector(15 downto 0);
        R_DATA          : out    vl_logic_vector(15 downto 0);
        ra              : out    vl_logic_vector(15 downto 0);
        rb              : out    vl_logic_vector(15 downto 0);
        temp            : out    vl_logic_vector(47 downto 0)
    );
end MyCPU;
