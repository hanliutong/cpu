library verilog;
use verilog.vl_types.all;
entity MY_REG_vlg_vec_tst is
end MY_REG_vlg_vec_tst;
