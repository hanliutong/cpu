library verilog;
use verilog.vl_types.all;
entity MyCPU_vlg_vec_tst is
end MyCPU_vlg_vec_tst;
