library verilog;
use verilog.vl_types.all;
entity registers_vlg_vec_tst is
end registers_vlg_vec_tst;
