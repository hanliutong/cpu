library verilog;
use verilog.vl_types.all;
entity CPU_Cycle_vlg_vec_tst is
end CPU_Cycle_vlg_vec_tst;
