library verilog;
use verilog.vl_types.all;
entity Memory_vlg_vec_tst is
end Memory_vlg_vec_tst;
