module tr(ADDC,SUBC,ANDC,ORC,XORC,NOTC,INCAC,DECAC,S3,S2,S1,S0,M,CN0);
input ADDC,SUBC,ANDC,ORC,XORC,NOTC,INCAC,DECAC;
output reg S3,S2,S1,S0,M,CN0;
always @ (ADDC or SUBC or ANDC or ORC or XORC or NOTC or INCAC or DECAC)
begin
	case({ADDC,SUBC,ANDC,ORC,XORC,NOTC,INCAC,DECAC})
		8'b00000001:{S3,S2,S1,S0,M,CN0} = 6'b111101;
		8'b00000010:{S3,S2,S1,S0,M,CN0} = 6'b000000;
		8'b00000100:{S3,S2,S1,S0,M,CN0} = 6'b00001x;
		8'b00001000:{S3,S2,S1,S0,M,CN0} = 6'b01101x;
		8'b00010000:{S3,S2,S1,S0,M,CN0} = 6'b11101x;
		8'b00100000:{S3,S2,S1,S0,M,CN0} = 6'b10111x;
		8'b01000000:{S3,S2,S1,S0,M,CN0} = 6'b011000;
		8'b10000000:{S3,S2,S1,S0,M,CN0} = 6'b100101;
		default: {S3,S2,S1,S0,M,CN0} = 6'b00111x;
	endcase
end
endmodule
