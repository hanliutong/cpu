library verilog;
use verilog.vl_types.all;
entity CLK_maker_vlg_vec_tst is
end CLK_maker_vlg_vec_tst;
