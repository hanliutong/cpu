library verilog;
use verilog.vl_types.all;
entity MyCPU_vlg_check_tst is
    port(
        A_plus          : in     vl_logic_vector(15 downto 0);
        ABUS            : in     vl_logic_vector(15 downto 0);
        ADDC            : in     vl_logic;
        ALU_IBUS        : in     vl_logic;
        BUS_MDR         : in     vl_logic;
        CLK             : in     vl_logic;
        cnt             : in     vl_logic_vector(3 downto 0);
        DBUS            : in     vl_logic_vector(15 downto 0);
        DECAC           : in     vl_logic;
        DST             : in     vl_logic;
        EXC             : in     vl_logic;
        FI              : in     vl_logic;
        I_DBUS          : in     vl_logic;
        IBUS            : in     vl_logic_vector(15 downto 0);
        IBUS_IR         : in     vl_logic;
        IBUS_MAR        : in     vl_logic;
        IBUS_PC         : in     vl_logic;
        IBUS_RA         : in     vl_logic;
        IBUS_RB         : in     vl_logic;
        IBUS_RBL        : in     vl_logic;
        IBUS_SR         : in     vl_logic;
        INCAC           : in     vl_logic;
        INT             : in     vl_logic;
        jieguo          : in     vl_logic_vector(15 downto 0);
        M_clk           : in     vl_logic;
        MAR_ABUS        : in     vl_logic;
        MAR_IBUS        : in     vl_logic;
        MDR_DBUS        : in     vl_logic;
        MDR_IBUS        : in     vl_logic;
        MRD             : in     vl_logic;
        MWR             : in     vl_logic;
        OpCode          : in     vl_logic_vector(5 downto 0);
        PC_IBUS         : in     vl_logic;
        PCplus1         : in     vl_logic;
        R               : in     vl_logic_vector(15 downto 0);
        R_DATA          : in     vl_logic_vector(15 downto 0);
        R_IBUS          : in     vl_logic;
        ra              : in     vl_logic_vector(15 downto 0);
        rb              : in     vl_logic_vector(15 downto 0);
        RBL_IBUS        : in     vl_logic;
        RE              : in     vl_logic;
        setTp1          : in     vl_logic;
        SR_IBUS         : in     vl_logic;
        SRC             : in     vl_logic;
        SUBC            : in     vl_logic;
        T               : in     vl_logic_vector(7 downto 0);
        temp            : in     vl_logic_vector(47 downto 0);
        W_B             : in     vl_logic;
        WE              : in     vl_logic;
        zero_PC         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MyCPU_vlg_check_tst;
