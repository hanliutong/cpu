module REGW2R(_reg,w,R);
input [2:0]_reg;
input w;
output reg [15:0]R;

always @ (_reg or w)
begin
	case({_reg,w})
	4'b000_0:R=16'b1000000000000000;
	4'b000_1:R=16'b0100000000000000;
	4'b001_0:R=16'b0010000000000000;
	4'b001_1:R=16'b0001000000000000;
	4'b010_0:R=16'b0000100000000000;
	4'b010_1:R=16'b0000010000000000;
	4'b011_0:R=16'b0000001000000000;
	4'b011_1:R=16'b0000000100000000;
	4'b100_0:R=16'b0000000010000000;
	4'b100_1:R=16'b0000000001000000;
	4'b101_0:R=16'b0000000000100000;
	4'b101_1:R=16'b0000000000010000;
	4'b110_0:R=16'b0000000000001000;
	4'b110_1:R=16'b0000000000000100;
	4'b111_0:R=16'b0000000000000010;
	4'b111_1:R=16'b0000000000000001;
	default:R=16'b000000000000000;
	endcase
end
endmodule

 