library verilog;
use verilog.vl_types.all;
entity CU_Timer_vlg_vec_tst is
end CU_Timer_vlg_vec_tst;
